package router_test_pkg;

import uvm_pkg::*;

`include "uvm_macros.svh"
`include "tb_defs.sv"
`include "source_xtn.sv"
`include "source_agent_config.sv"
`include "destination_agent_config.sv"
`include "router_env_config.sv"
`include "source_driver.sv"
`include "source_monitor.sv"
`include "source_sequencer.sv"
`include "source_agent.sv"
`include "source_agt_top.sv"
`include "source_seqs.sv"


`include "destination_xtn.sv"
`include "destination_monitor.sv"
`include "destination_sequencer.sv"
`include "destination_seqs.sv"
`include "destination_driver.sv"
`include "destination_agent.sv"
`include "destination_agt_top.sv"

`include "router_virtual_sequencer.sv"
`include "router_virtual_seqs.sv"
`include "router_scoreboard.sv"

`include "router_tb.sv"


`include "router_vtest_lib.sv"
endpackage
